module soupbintcp3{

}{
	input clk,
	input nreset
}

endmodule; 
